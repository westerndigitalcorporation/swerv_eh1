// NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE
// This is an automatically generated file by joseph.rahmeh on Tue Jun  4 07:50:46 PDT 2019
//
// cmd:    swerv -snapshot=default -ahb_lite 
//

`include "common_defines.vh"
`undef ASSERT_ON
`undef TEC_RV_ICG
`define TEC_RV_ICG CKLNQD12BWP35P140
`define PHYSICAL 1
